//A function to check if the CRC is correct according to 6

