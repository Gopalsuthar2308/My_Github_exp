//5.1 write a class as packet which has function which will give count of how many times packet is generated.
//5.2 modify function in Q1 with automatic function and what will be the difference between the outpug.
